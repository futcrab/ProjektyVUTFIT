library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
library work;

entity MEMORY is
Port ( INDEX 		: in INTEGER;
       COL_VALUE  : out STD_LOGIC_VECTOR(7 downto 0)); 
end MEMORY;

architecture Behavioral of MEMORY is
-- smile face bitmap   00000000 00000000 00011000 00100000 01000000 01001110 11000000 11000000 11000000 11000000 01001110 01000000 00100000 00011000 00000000 00000000
--							  00000000 00000010 00000110 00010110 00001110 00101110 11111011 00000010 11111011 00101110 00001110 00010110 00000110 00000010 00000000 00000000
--							  00000000 00000000 10000000 11000000 11111100 00110010 00010001 00010101 00010001 00110010 11111100 11000000 10000000 00000000 00000000 00000000
--							  00000000 00000000 00000000 00010000 00101000 00101000 01000100 10000010 11101110 00101000 00101000 00111100 00000000 00000000 00000000 00000000
--							  00000000 00000000 00000000 00111100 01000010 10111101 10000101 10111101 10000101 10111101 01000010 00111100 00000000 00000000 00000000 00000000

type DATA is array (0 to 63) of std_logic_vector(7 downto 0);

		                
constant MEMORY: DATA := 
(
		"00000000", "00000010", "00000110", "00010110", "00001110", "00101110", "11111011", "00000010", "11111011", "00101110", "00001110", "00010110","00000110", "00000010", "00000000", "00000000",
		"00000000", "00000000", "10000000", "11000000", "11111100", "00110010", "00010001", "00010101", "00010001", "00110010", "11111100", "11000000", "10000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00010000", "00101000", "00101000", "01000100", "10000010", "11101110", "00101000", "00101000", "00111100", "00000000", "00000000", "00000000", "00000000",
	   "00000000", "00000000", "00000000", "00111100", "01000010", "10111101", "10100001", "10111101", "10100001", "10111101", "01000010", "00111100", "00000000", "00000000", "00000000", "00000000"
);

begin
	COL_VALUE <= MEMORY(INDEX);
end Behavioral;