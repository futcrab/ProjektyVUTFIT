LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.effects_pack.ALL;
LIBRARY work;

ENTITY stlpec IS
	PORT (
		CLK : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		STATE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		INIT_STATE : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		NEIGH_LEFT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		NEIGH_RIGHT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		DIRECTION : IN DIRECTION_T;
		EN : IN STD_LOGIC);
END stlpec;

ARCHITECTURE Behavioral OF stlpec IS

BEGIN
	PROCESS (CLK)
	BEGIN
		IF rising_edge(CLK) THEN
			IF RESET = '1' THEN
				STATE <= INIT_STATE;
			ELSIF EN = '1' THEN
				IF DIRECTION = DIR_RIGHT THEN
					STATE <= NEIGH_RIGHT;
				ELSIF DIRECTION = DIR_LEFT THEN
					STATE <= NEIGH_LEFT;
				ELSIF DIRECTION = DIR_TOP THEN
					STATE <= INIT_STATE(0) & INIT_STATE(7 DOWNTO 1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
END Behavioral;